.title KiCad schematic
.include "/usr/share/kicad/models/1N5818.mod"
.include "/usr/share/kicad/models/TL074.mod"
D2 GNDPWR -v 1N5818
C7 +v GNDPWR 0.1uf
C2 GNDPWR -v 10uf
C8 -v GNDPWR 0.1uf
C1 +v GNDPWR 10uf
R12 Output12 Net-_R12-Pad2_ 1k
D1 +v GNDPWR 1N5818
C6 -v GNDPWR 0.1uf
C5 +v GNDPWR 0.1uf
C3 +v GNDPWR 0.1uf
C4 -v GNDPWR 0.1uf
R13 Output11 Net-_R12-Pad2_ 1k
R14 Output10 Net-_R14-Pad2_ 1k
R11 Output9 Net-_R11-Pad2_ 1k
XU3 Net-_R11-Pad2_ Net-_R11-Pad2_ InputBus3 +v InputBus4 Net-_R14-Pad2_ Net-_R14-Pad2_ Net-_U3-Pad8_ Net-_U3-Pad8_ InputBus4 -v InputBus4 Net-_R12-Pad2_ Net-_R12-Pad2_ TL074
R4 Output4 Net-_R4-Pad2_ 1k
R3 Output3 Net-_R3-Pad2_ 1k
R1 Output1 Net-_R1-Pad2_ 1k
R2 Output2 Net-_R2-Pad2_ 1k
Vin1 InputBus1 GNDPWR dc 1 sin(0 3 1k 0 0 0)
XU1 Net-_R1-Pad2_ Net-_R1-Pad2_ InputBus1 +v InputBus1 Net-_R2-Pad2_ Net-_R2-Pad2_ Net-_R3-Pad2_ Net-_R3-Pad2_ InputBus1 -v InputBus2 Net-_R4-Pad2_ Net-_R4-Pad2_ TL074
XU2 Net-_R5-Pad2_ Net-_R5-Pad2_ InputBus2 +v InputBus2 Net-_R6-Pad2_ Net-_R6-Pad2_ Net-_R7-Pad2_ Net-_R7-Pad2_ InputBus3 -v InputBus3 Net-_R8-Pad2_ Net-_R8-Pad2_ TL074
R6 Output6 Net-_R6-Pad2_ 1k
R5 Output5 Net-_R5-Pad2_ 1k
R7 Output7 Net-_R7-Pad2_ 1k
R8 Output8 Net-_R8-Pad2_ 1k
.op
.control
.options rshunt=100M gmin=10n
tran 99.999us 1.005s 1s
set color0=rgb:f/f/f
set color1=rgb:0/0/0
set color2=rgb:0/0/f
set color3=rgb:f/f/0
set color4=rgb:0/f/f
set color5=rgb:f/0/f
set color6=rgb:5/0/0
hardcopy BufferedMultiple.ps V(InputBus1) V(Output1) V(Output2) V(output3) V(Output4)
.endc
.end
